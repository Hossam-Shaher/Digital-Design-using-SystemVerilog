module buffer (
  input [15:0] I,		//input wire logic [15:0]
  output [15:0] O		//output wire logic [15:0]
);
  
  assign O = I;
  
endmodule: buffer